module pmod_ad1_wrapper (
  input CLK_i,
  output AD7476_CS_o,
  output AD7476_SCLK_o,
  input AD7476_SDATA0_i,
  input AD7476_SDATA1_i,
  output [15:0] ADC_DATA0_o,
  output [15:0] ADC_DATA1_o,
  output ADC_VALID_o,
  //AXI4-Stream Interface
  output [15:0] M_AXIS_TDATA,
  output [1:0] M_AXIS_TKEEP,
  output M_AXIS_TLAST,
  input M_AXIS_TREADY,
  output M_AXIS_TVALID,
  //AXI4-Lite Interface
  input AXI_ACLK_i,
  input AXI_ARESETN_i,
  input [31:0] S_AXI_ARADDR,
  output S_AXI_ARREADY,
  input S_AXI_ARVALID,
  input [31:0] S_AXI_AWADDR,
  output S_AXI_AWREADY,
  input S_AXI_AWVALID,
  input S_AXI_BREADY,
  output [1:0] S_AXI_BRESP,
  output S_AXI_BVALID,
  output [31:0] S_AXI_RDATA,
  input S_AXI_RREADY,
  output [1:0] S_AXI_RRESP,
  output S_AXI_RVALID,
  input [31:0] S_AXI_WDATA,
  output S_AXI_WREADY,
  input [3:0] S_AXI_WSTRB,
  input S_AXI_WVALID
);

pmod_ad1 pmod_ad1_inst (
  .CLK_i           (CLK_i),
  .AD7476_CS_o     (AD7476_CS_o),
  .AD7476_SCLK_o   (AD7476_SCLK_o),
  .AD7476_SDATA0_i (AD7476_SDATA0_i),
  .AD7476_SDATA1_i (AD7476_SDATA1_i),
  .ADC_DATA0_o     (ADC_DATA0_o),
  .ADC_DATA1_o     (ADC_DATA1_o),
  .ADC_VALID_o     (ADC_VALID_o),
  //AXI4-Stream Interface
  .AXIS_TDATA_o    (M_AXIS_TDATA),
  .AXIS_TKEEP_o    (M_AXIS_TKEEP),
  .AXIS_TLAST_o    (M_AXIS_TLAST),
  .AXIS_TREADY_i   (M_AXIS_TREADY),
  .AXIS_TVALID_o   (M_AXIS_TVALID),
  //AXI4-Lite Interface
  .AXI_ACLK_i      (AXI_ACLK_i),
  .AXI_ARESETN_i   (AXI_ARESETN_i),
  .AXI_ARADDR_i    (S_AXI_ARADDR),
  .AXI_ARREADY_o   (S_AXI_ARREADY),
  .AXI_ARVALID_i   (S_AXI_ARVALID),
  .AXI_AWADDR_i    (S_AXI_AWADDR),
  .AXI_AWREADY_o   (S_AXI_AWREADY),
  .AXI_AWVALID_i   (S_AXI_AWVALID),
  .AXI_BREADY_i    (S_AXI_BREADY),
  .AXI_BRESP_o     (S_AXI_BRESP),
  .AXI_BVALID_o    (S_AXI_BVALID),
  .AXI_RDATA_o     (S_AXI_RDATA),
  .AXI_RREADY_i    (S_AXI_RREADY),
  .AXI_RRESP_o     (S_AXI_RRESP),
  .AXI_RVALID_o    (S_AXI_RVALID),
  .AXI_WDATA_i     (S_AXI_WDATA),
  .AXI_WREADY_o    (S_AXI_WREADY),
  .AXI_WSTRB_i     (S_AXI_WSTRB),
  .AXI_WVALID_i    (S_AXI_WVALID)
);

endmodule
